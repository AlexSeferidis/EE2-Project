module single_engine (
    input logic clk,
    input logic reset,
    input logic [31:0] iterations_max,
    input logic signed [fp_bits - 1:0] x0,
    input logic signed [fp_bits - 1:0] y0,

    output logic finished,
    output logic [31:0] iterations
  );









endmodule
